module const128 (
output [31:0] result
);
assign result = 32'b01000011000000000000000000000000;
endmodule